library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FlipFlopD_tb is
end FlipFlopD_tb;

architecture teste of FlipFlopD_tb is

   component FlipFlopD is
	port( clock: in std_logic;
		  D: in std_logic;
		  reset: in std_logic;
	      Q : inout std_logic :='0';
			Qi: inout std_logic :='0'
	    );
end component;

signal clock, D, reset : std_logic;
signal Q, Qi : std_logic := '0';
signal   running		 : bit;
 
begin

flip_flop : FlipFlopD port map (clock => clock, D => D, reset => reset, Q =>Q, Qi=>Qi);

running <= '1', '0' after 50 ns; 

clock <= not clock after 3 ns when running = '1' else '0';
D <= '0', '1' after 2 ns, '0' after 5 ns, '1' after 11 ns, '0' after 17 ns, '1' after 22 ns, '0' after 25 ns, '1' after 30 ns, '0' after 35 ns;
reset <= '0';

end teste;